module Hazard_Detection_Sim;
    
endmodule